`default_nettype none


module waveshaper(
    //inputs
    //outputs
);

//internal signals

//your code here

endmodule


module sequential_div(
    //inputs
    //outputs
);

//internal signals

//your code here

endmodule
