`default_nettype none


module sample_rate_clkdiv(
    //inputs
    //outputs
);

//internal signals

//your code here

endmodule
```