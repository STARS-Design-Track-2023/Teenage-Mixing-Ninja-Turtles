`default_nettype none


module pwm(
    //inputs
    //outputs
);

//internal signals

//your code here

endmodule
```