
module oscillator(
    //inputs
    //outputs
);

//internal signals

// your code goes here

endmodule
```