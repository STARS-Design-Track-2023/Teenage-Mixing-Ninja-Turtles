`default_nettype none


module keypad(
    //inputs
    //outputs
);

//internal signals

//your code here

endmodule
```