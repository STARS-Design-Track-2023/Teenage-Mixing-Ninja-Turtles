`default_nettype none


module signal_mixr(
    //inputs
    //outputs
);

//internal signals

//your code here

endmodule
